/////////////////////////////////////////////////////////////////////////
//                                                                     //
//                                                                     //
//   Modulename :  testbench.v                                         //
//                                                                     //
//  Description :  Testbench module for the verisimple pipeline;       //
//                                                                     //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

`timescale 1ns/100ps
extern void print_header(string str);
extern void print_cycles();
extern void print_stage(string div, int inst, int npc, int valid_inst);
extern void print_reg(int wb_reg_wr_data_out_hi, int wb_reg_wr_data_out_lo,
                      int wb_reg_wr_idx_out, int wb_reg_wr_en_out);
extern void print_membus(int proc2mem_command, int mem2proc_response,
                         int proc2mem_addr_hi, int proc2mem_addr_lo,
                         int proc2mem_data_hi, int proc2mem_data_lo);
extern void print_close();
extern void print_cycles_same();

module testbench;

  // variables used in the testbench
  logic        clock;
  logic        reset;
  logic [31:0] clock_count;
  logic [31:0] instr_count;
  int          wb_fileno;

  logic [1:0]  proc2mem_command;
  logic [63:0] proc2mem_addr;
  logic [63:0] proc2mem_data;
  logic  [3:0] mem2proc_response;
  logic [63:0] mem2proc_data;
  logic  [3:0] mem2proc_tag;

  logic  [3:0] pipeline_completed_insts_0,pipeline_completed_insts_1;
  ERROR_CODE  pipeline_error_status;
  logic  [$clog2(`N_ENTRY_ROB+33)-1:0] pipeline_commit_wr_idx_0, pipeline_commit_wr_idx_1;
  logic [63:0] pipeline_commit_wr_data_0, pipeline_commit_wr_data_1;
  logic        pipeline_commit_wr_en_0, pipeline_commit_wr_en_1;
  logic [63:0] pipeline_commit_NPC_0, pipeline_commit_NPC_1;


  logic [63:0] if_NPC_out_0;
  logic [31:0] if_IR_out_0;
  logic        if_valid_inst_out_0;
  logic [63:0] if_NPC_out_1;
  logic [31:0] if_IR_out_1;
  logic        if_valid_inst_out_1;
  logic [63:0] if_id_NPC_0;
  logic [31:0] if_id_IR_0;
  logic        if_id_valid_inst_0;
  logic [63:0] if_id_NPC_1;
  logic [31:0] if_id_IR_1;
  logic        if_id_valid_inst_1;
  logic [63:0] id_ex_NPC_0;
  logic [31:0] id_ex_IR_0;
  logic        id_ex_valid_inst_0;
  logic [63:0] id_ex_NPC_1;
  logic [31:0] id_ex_IR_1;
  logic        id_ex_valid_inst_1;
  logic [63:0] ex_mem_NPC_0;
  logic [31:0] ex_mem_IR_0;
  logic        ex_mem_valid_inst_0;
  logic [63:0] ex_mem_NPC_1;
  logic [31:0] ex_mem_IR_1;
  logic        ex_mem_valid_inst_1;
  logic [63:0] mem_wb_NPC_0;
  logic [31:0] mem_wb_IR_0;
  logic        mem_wb_valid_inst_0;
  logic [63:0] mem_wb_NPC_1;
  logic [31:0] mem_wb_IR_1;
  logic        mem_wb_valid_inst_1;

  logic valid_wb_0;
  logic valid_wb_1; //valid bit

// add
logic 	[31:0][63:0] test_rf_value;
logic	[4:0] wr_idx_0_out;
logic	[4:0] wr_idx_1_out;
logic	[63:0] wr_value_0_out;
logic	[63:0] wr_value_1_out;
logic	retire_valid_0_out;
logic	retire_valid_1_out;
logic	[63:0] retire_NPC_0_out;
logic	[63:0] retire_NPC_1_out;

logic [63:0] ROB_rt_NPC_out_0;
logic [63:0] ROB_rt_NPC_out_1;
logic [31:0] ROB_rt_IR_out_0;
logic [31:0] ROB_rt_IR_out_1;


logic [31:0] [$clog2(`N_ENTRY_ROB+33)-1:0] rt_tag_out;
logic [`N_ENTRY_ROB+32:0][63:0] rf_value_out;
logic free_PR_1;
logic free_PR_0;
logic [4:0] wr_idx_0;
logic [4:0] wr_idx_1;
logic [$clog2(`N_ENTRY_ROB+33)-1:0] rt_Tnew_out_0;
logic [$clog2(`N_ENTRY_ROB+33)-1:0] rt_Tnew_out_1;
logic [$clog2(`N_ENTRY_ROB+33)-1:0] rt_Told_out_0;
logic [$clog2(`N_ENTRY_ROB+33)-1:0] rt_Told_out_1;

logic is_0_br;
logic recovery_request;
logic [$clog2(`N_ENTRY_ROB)-1:0] recovery_tail;
logic [$clog2(`N_ENTRY_ROB+33)-1:0] free_list_in_0;
logic [$clog2(`N_ENTRY_ROB+33)-1:0] free_list_in_1;
logic [$clog2(`N_ENTRY_ROB+33)-1:0] CDB_in_0; 
logic [$clog2(`N_ENTRY_ROB+33)-1:0] CDB_in_1; 
logic [$clog2(`N_ENTRY_ROB+33)-1:0] T_old_0;
logic [$clog2(`N_ENTRY_ROB+33)-1:0] T_old_1;
logic fetch_PR_0;
logic fetch_PR_1;
logic id_halt_out_0;
logic id_halt_out_1;
logic id_wr_mem_out_0;
logic id_wr_mem_out_1;




  // Instantiate the Pipeline
  pipeline pipeline_0 (
    //ah hahahahahaha
	.rf_value_out(rf_value_out),
	.free_PR_1(free_PR_1),
	.free_PR_0(free_PR_0),
  .rt_Told_out_0(rt_Told_out_0),
  .rt_Told_out_1(rt_Told_out_1),
  .rt_Tnew_out_0(rt_Tnew_out_0),
  .rt_Tnew_out_1(rt_Tnew_out_1),
	.is_0_br(is_0_br),
	.recovery_request(recovery_request),
	.recovery_tail(recovery_tail),
	.free_list_in_0(free_list_in_0),
	.free_list_in_1(free_list_in_1),
	.CDB_in_0(CDB_in_0),
	.CDB_in_1(CDB_in_1),
	.T_old_0(T_old_0),
	.T_old_1(T_old_1),
	.fetch_PR_0(fetch_PR_0),
	.fetch_PR_1(fetch_PR_1),
	.id_halt_out_0(id_halt_out_0),
	.id_halt_out_1(id_halt_out_1),
	.id_wr_mem_out_0(id_wr_mem_out_0),
	.id_wr_mem_out_1(id_wr_mem_out_1),

    // Inputs
    .clock             (clock),
    .reset             (reset),
    .mem2proc_response (mem2proc_response),
    .mem2proc_data     (mem2proc_data),
    .mem2proc_tag      (mem2proc_tag),
    //

    .valid_wb_0(valid_wb_0),
    .valid_wb_1(valid_wb_1), //valid bit
    // Outputs

    .proc2mem_command  (proc2mem_command),
    .proc2mem_addr     (proc2mem_addr),
    .proc2mem_data     (proc2mem_data),

    .pipeline_completed_insts_0(pipeline_completed_insts_0),
    .pipeline_error_status(pipeline_error_status),
    .pipeline_commit_wr_data_0(pipeline_commit_wr_data_0),
    .pipeline_commit_wr_idx_0(pipeline_commit_wr_idx_0),
    .pipeline_commit_wr_en_0(pipeline_commit_wr_en_0),
    .pipeline_commit_NPC_0(pipeline_commit_NPC_0),

    .if_NPC_out_0(if_NPC_out_0),
    .if_IR_out_0(if_IR_out_0),
    .if_valid_inst_out_0(if_valid_inst_out_0),
    .if_id_NPC_0(if_id_NPC_0),
    .if_id_IR_0(if_id_IR_0),
    .if_id_valid_inst_0(if_id_valid_inst_0),
    .id_ex_NPC_0(id_ex_NPC_0),
    .id_ex_IR_0(id_ex_IR_0),
    .id_ex_valid_inst_0(id_ex_valid_inst_0),
    .ex_mem_NPC_0(ex_mem_NPC_0),
    .ex_mem_IR_0(ex_mem_IR_0),
    .ex_mem_valid_inst_0(ex_mem_valid_inst_0),

    .pipeline_completed_insts_1(pipeline_completed_insts_1),
    .pipeline_commit_wr_data_1(pipeline_commit_wr_data_1),
    .pipeline_commit_wr_idx_1(pipeline_commit_wr_idx_1),
    .pipeline_commit_wr_en_1(pipeline_commit_wr_en_1),
    .pipeline_commit_NPC_1(pipeline_commit_NPC_1),

    .if_NPC_out_1(if_NPC_out_1),
    .if_IR_out_1(if_IR_out_1),
    .if_valid_inst_out_1(if_valid_inst_out_1),
    .if_id_NPC_1(if_id_NPC_1),
    .if_id_IR_1(if_id_IR_1),
    .if_id_valid_inst_1(if_id_valid_inst_1),
    .id_ex_NPC_1(id_ex_NPC_1),
    .id_ex_IR_1(id_ex_IR_1),
    .id_ex_valid_inst_1(id_ex_valid_inst_1),
    .ex_mem_NPC_1(ex_mem_NPC_1),
    .ex_mem_IR_1(ex_mem_IR_1),
    .ex_mem_valid_inst_1(ex_mem_valid_inst_1)

    //For DEBUG

  );

  ArchMap ArchMap_0(
    .clock(clock),
    .reset(reset),
    .valid_0(free_PR_0),
    .valid_1(free_PR_1),
    .Told_out_0(rt_Told_out_0), 
    .Told_out_1(rt_Told_out_1),
    .Tnew_out_0(rt_Tnew_out_0),
    .Tnew_out_1(rt_Tnew_out_1),

    .tag(rt_tag_out),   //modified for test
    .wr_idx_0(wr_idx_0),  //modified for test
    .wr_idx_1(wr_idx_1)   //modified for test
  );

  test_reg test_reg0(
	.clk(clock),
	.rst(reset),
	.tag(rt_tag_out),
	.value_RF(rf_value_out),
	.valid_1(free_PR_1),
	.valid_0(free_PR_0),
	.wr_idx_0(wr_idx_0),
	.wr_idx_1(wr_idx_1),
	.Tnew_out_0(rt_Tnew_out_0),
	.Tnew_out_1(rt_Tnew_out_1),
	.retire_NPC_0_in(ROB_rt_NPC_out_0),
	.retire_NPC_1_in(ROB_rt_NPC_out_1),

	.test_rf_value(test_rf_value),
	.wr_idx_0_out(wr_idx_0_out),
	.wr_idx_1_out(wr_idx_1_out),
	.wr_value_0_out(wr_value_0_out),
	.wr_value_1_out(wr_value_1_out),

	.retire_valid_0_out(retire_valid_0_out),
	.retire_valid_1_out(retire_valid_1_out),
	.retire_NPC_0_out(retire_NPC_0_out),
	.retire_NPC_1_out(retire_NPC_1_out)
  ); 


 ROB_test ROB_test (
    .clock(clock),
    .reset(reset),
    .is_0_br(is_0_br),
    .recovery_br(recovery_request),///////from EX-mem stage
    .recovery_tail(recovery_tail),
    .freelist_0(free_list_in_0), .freelist_1(free_list_in_1),
    .CDB_in_0(CDB_in_0), .CDB_in_1(CDB_in_1),
    .map_table_Told_in_0(T_old_0),
    .map_table_Told_in_1(T_old_1),
    .fetch_PR_0(fetch_PR_0),
    .fetch_PR_1(fetch_PR_1),
    .ROB_halt_in_0(id_halt_out_0),
    .ROB_halt_in_1(id_halt_out_1),
    .is_0_st(id_wr_mem_out_0),
    .is_1_st(id_wr_mem_out_1),
    .if_id_NPC_0(if_id_NPC_0), .if_id_NPC_1(if_id_NPC_1),
	.if_id_IR_0(if_id_IR_0), .if_id_IR_1(if_id_IR_1),

	// Output
    .ROB_rt_NPC_out_0(ROB_rt_NPC_out_0),
    .ROB_rt_NPC_out_1(ROB_rt_NPC_out_1),
    .ROB_rt_IR_out_0(ROB_rt_IR_out_0),
    .ROB_rt_IR_out_1(ROB_rt_IR_out_1)
  );




  // Instantiate the Data Memory
  mem memory (
    // Inputs
    .clk               (clock),
    .proc2mem_command  (proc2mem_command),
    .proc2mem_addr     (proc2mem_addr),
    .proc2mem_data     (proc2mem_data),

    // Outputs

    .mem2proc_response (mem2proc_response),
    .mem2proc_data     (mem2proc_data),
    .mem2proc_tag      (mem2proc_tag)
  );

  parameter REG_IDX_0_FILL = 32 - $clog2(`N_ENTRY_ROB+33);
  // Generate System Clock
  always begin
    #(`VERILOG_CLOCK_PERIOD/2.0);
    clock = ~clock;
  end

  // Task to display # of elapsed clock edges
  task show_clk_count;
    real cpi;

    begin
      cpi = (clock_count + 1.0) / instr_count;
      $display("@@  %0d cycles / %0d instrs = %f CPI\n@@",
                clock_count+1, instr_count, cpi);
      $display("@@  %4.2f ns total time to execute\n@@\n",
                clock_count*`VIRTUAL_CLOCK_PERIOD);
    end
  endtask  // task show_clk_count

  // Show contents of a range of Unified Memory, in both hex and decimal
  task show_mem_with_decimal;
    input [31:0] start_addr;
    input [31:0] end_addr;
    int showing_data;
    begin
      $display("@@@");
      showing_data=0;
      for(int k=start_addr;k<=end_addr; k=k+1)
        if (memory.unified_memory[k] != 0) begin
          $display("@@@ mem[%5d] = %x : %0d", k*8, memory.unified_memory[k], 
                                                    memory.unified_memory[k]);
          showing_data=1;
        end else if(showing_data!=0) begin
          $display("@@@");
          showing_data=0;
        end
      $display("@@@");
    end
  endtask  // task show_mem_with_decimal

  initial begin
  
    clock = 1'b0;
    reset = 1'b0;

    // Pulse the reset signal
    $display("@@\n@@\n@@  %t  Asserting System reset......", $realtime);
    reset = 1'b1;
    @(posedge clock);
    @(posedge clock);

    $readmemh("program.mem", memory.unified_memory);

    @(posedge clock);
    @(posedge clock);
    `SD;
    // This reset is at an odd time to avoid the pos & neg clock edges

    reset = 1'b0;
    $display("@@  %t  Deasserting System reset......\n@@\n@@", $realtime);

    wb_fileno = $fopen("writeback.out");
    
    //Open header AFTER throwing the reset otherwise the reset state is displayed
    print_header("                                                                            D-MEM Bus &\n");
    print_header("Cycle:      IF      |     ID      |     EX      |     CPL     |     RT      Reg Result");
  end


  // Count the number of posedges and number of instructions completed
  // till simulation ends
  always @(posedge clock) begin
    if(reset) begin
      clock_count <= `SD 0;
      instr_count <= `SD 0;
    end else begin
      clock_count <= `SD (clock_count + 1);
      //instr_count <= `SD (instr_count + pipeline_completed_insts_0 + pipeline_completed_insts_0);
      instr_count <= `SD (instr_count + valid_wb_0 + valid_wb_1);
    end
  end  


  always @(negedge clock) begin
    if(reset)
      $display("@@\n@@  %t : System STILL at reset, can't show anything\n@@",
               $realtime);
    else begin
      `SD;
      `SD;
      
       // print the piepline stuff via c code to the pipeline.out
       print_cycles();
       print_stage(" ", if_IR_out_0, if_NPC_out_0[31:0], {31'b0,if_valid_inst_out_0});
       print_stage("|", if_id_IR_0, if_id_NPC_0[31:0], {31'b0,if_id_valid_inst_0});
       print_stage("|", id_ex_IR_0, id_ex_NPC_0[31:0], {31'b0,id_ex_valid_inst_0});
       print_stage("|", ex_mem_IR_0, ex_mem_NPC_0[31:0], {31'b0,ex_mem_valid_inst_0});
       print_stage("|", ROB_rt_IR_out_0, ROB_rt_NPC_out_0[31:0], {31'b0,valid_wb_0});
       print_reg(pipeline_commit_wr_data_0[63:32], pipeline_commit_wr_data_0[31:0],
                 {{REG_IDX_0_FILL{1'b0}},pipeline_commit_wr_idx_0}, {31'b0,pipeline_commit_wr_en_0});
       // TO DO
       print_membus({30'b0,proc2mem_command}, {28'b0,mem2proc_response},
                    proc2mem_addr[63:32], proc2mem_addr[31:0],
                    proc2mem_data[63:32], proc2mem_data[31:0]);
       print_cycles_same();
       print_stage(" ", if_IR_out_1, if_NPC_out_1[31:0], {31'b0,if_valid_inst_out_1});
       print_stage("|", if_id_IR_1, if_id_NPC_1[31:0], {31'b0,if_id_valid_inst_1});
       print_stage("|", id_ex_IR_1, id_ex_NPC_1[31:0], {31'b0,id_ex_valid_inst_1});
       print_stage("|", ex_mem_IR_1, ex_mem_NPC_1[31:0], {31'b0,ex_mem_valid_inst_1});
       print_stage("|", ROB_rt_IR_out_1, ROB_rt_NPC_out_1[31:0], {31'b0,valid_wb_1});
       print_reg(pipeline_commit_wr_data_1[63:32], pipeline_commit_wr_data_1[31:0],
                 {{REG_IDX_0_FILL{1'b0}},pipeline_commit_wr_idx_1}, {31'b0,pipeline_commit_wr_en_1});
       // TO DO
       print_membus({30'b0,proc2mem_command}, {28'b0,mem2proc_response},
                    proc2mem_addr[63:32], proc2mem_addr[31:0],
                    proc2mem_data[63:32], proc2mem_data[31:0]);


      if(retire_valid_0_out) begin
        if (wr_idx_0_out != `ZERO_REG) begin
          $fdisplay(wb_fileno, "PC=%x, REG[%d]=%x",
                    retire_NPC_0_out-4,
                    wr_idx_0_out,
                    wr_value_0_out);
        end else begin
          $fdisplay(wb_fileno, "PC=%x, ---",
                    retire_NPC_0_out-4);
        end
      end

      if(retire_valid_1_out) begin
        if (wr_idx_1_out != `ZERO_REG) begin
          $fdisplay(wb_fileno, "PC=%x, REG[%d]=%x",
                     retire_NPC_1_out-4,
                     wr_idx_1_out,
                     wr_value_1_out);
        end else begin
          $fdisplay(wb_fileno, "PC=%x, ---",
                     retire_NPC_1_out-4);
        end
      end

      // deal with any halting conditions
      if(pipeline_error_status != NO_ERROR) begin
        $display("@@@ Unified Memory contents hex on left, decimal on right: ");
        show_mem_with_decimal(0,`MEM_64BIT_LINES - 1); 
          // 8Bytes per line, 16kB total

        $display("@@  %t : System halted\n@@", $realtime);

        case(pipeline_error_status)
          HALTED_ON_MEMORY_ERROR:  
              $display("@@@ System halted on memory error");
          HALTED_ON_HALT:          
              $display("@@@ System halted on HALT instruction");
          HALTED_ON_ILLEGAL:
              $display("@@@ System halted on illegal instruction");
          default: 
              $display("@@@ System halted on unknown error code %x",
                       pipeline_error_status);
        endcase
        $display("@@@\n@@");
        show_clk_count;
        print_close(); // close the pipe_print output file
        $fclose(wb_fileno);
        #100 $finish;
      end

    end  // if(reset)   
  end 

endmodule  // module testbench
